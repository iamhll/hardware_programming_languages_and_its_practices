// skip checkFileHeader
