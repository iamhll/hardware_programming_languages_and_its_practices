// CRC
`define CRC_NUMB_INP       'd1813
`define CRC_SIZE_POLY      'h12
`define CRC_DATA_POLY      'h1CF91
`define CRC_DATA_INIT      'h75C0A
`define CRC_DATA_XOROUT    'h77CEB
`define CRC_FLAG_REFIN     'h0
`define CRC_FLAG_REFOUT    'h1
