//------------------------------------------------------------------------------
  //
  //  Filename       : localparam_calc.vh
  //  Author         : Huang Leilei
  //  Status         : draft
  //  Created        : 2025-02-18
  //  Description    : [parameter] of [xkcalc]
  //
//------------------------------------------------------------------------------
